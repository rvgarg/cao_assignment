LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY 4bit_ripple_behavioural IS
    --  Port ( );
END 4bit_ripple_behavioural;

ARCHITECTURE Behavioral OF 4bit_ripple_behavioural IS

BEGIN
END Behavioral;